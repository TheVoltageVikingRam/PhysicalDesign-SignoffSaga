module tb;
reg [9:0] in;
reg [3:0] s;
wire y;

mux10 uut ( .in(in), .s(s), .y(y));

initial begin

in = 10'b1111111111; s = 4'd3; #10;
in = 10'b1111000111; s = 4'd2; #10;
in = 10'b1001111111; s = 4'd1; #10;
in = 10'b1111110111; s = 4'd4; #10;
in = 10'b1111011111; s = 4'd5; #10;
in = 10'b1110001111; s = 4'd6; #10;
in = 10'b1111100000; s = 4'd9; #10;
in = 10'b0000001111; s = 4'd3; #10;
in = 10'b1111111111; s = 4'd8; #10;
in = 10'b1111110000; s = 4'd7; #10;

$finish();


end
endmodule
